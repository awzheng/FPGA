module LogicalStep_Lab2_top
(
	input				rst_n,		//reset in
	input          clkin_50,	//clock in
	input		[7:0]	sw,
	input		[3:0]	pb_n,

	output	[7:0]	leds,
	output	[6:0]	seg7_data,
	output			seg7_char1,
	output			seg7_char2

);

//these are used as intermediate signals
	wire 	[3:0] hex_A, hex_B;
	wire	[6:0] seg7_A, seg7_B;
	wire 	[3:0] pb;

	
// wire assignments
	assign hex_A = sw[3:0];
	assign hex_B = sw[7:4];

	
//module instantiations are here
	SevenSegment u1 (
		.hex      (hex_A), 
		.sevenseg (seg7_A)
	);

	SevenSegment u2 (
		.hex      (hex_B), 
		.sevenseg (seg7_B)
	);

	segment7_mux u3 (
		.clk  (clkin_50),
		.din2 (seg7_A), 
		.din1 (seg7_B),
		.dout (seg7_data),
		.dig2 (seg7_char2), 
		.dig1 (seg7_char1)
	);
	
	pb_inverters u4 (
		.pbin  (pb_n),
		.pbout (pb)
	);
	
	mux_4bit_2_to_1 (
	
		.din_A (hex_A),
		.din_B (hex_B),
		.selector (pb[1:0]),
		.dout (leds[3:0])
	
	);
 
 
 
endmodule

	